-- Example VHDL source file
-- Example simulation VHDL file